////////////////////////////////////////////////////////
/////////////struct para los bits de paridad/////////////
////////////////////////////////////////////////////////
package hamming_pkg;
typedef struct packed {
  logic p1;
  logic p2;
  logic p3;
} hamming_parity_t;
endpackage
